/*------------------------------------------------------------------------------
 * File          : Pattern_Generator_sequencer.sv
 * Project       : RTL
 * Author        : epmkos
 * Creation date : Jul 30, 2024
 * Description   :
 *------------------------------------------------------------------------------*/

module Pattern_Generator_sequencer #() ();

endmodule