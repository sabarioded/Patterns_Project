/*------------------------------------------------------------------------------
 * File          : Pattern_Generator_driver.sv
 * Project       : RTL
 * Author        : epmkos
 * Creation date : Jul 30, 2024
 * Description   :
 *------------------------------------------------------------------------------*/

module Pattern_Generator_driver #() ();

endmodule